library verilog;
use verilog.vl_types.all;
entity combinacional_vlg_vec_tst is
end combinacional_vlg_vec_tst;
