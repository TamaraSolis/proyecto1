library verilog;
use verilog.vl_types.all;
entity negador_vlg_vec_tst is
end negador_vlg_vec_tst;
